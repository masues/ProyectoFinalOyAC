library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity u_control is
	Port( inst : in STD_LOGIC_VECTOR (15 downto 0);
			selregr : out STD_LOGIC_VECTOR (3 downto 0);
			sels1 : out STD_LOGIC;
			sr : out STD_LOGIC;
			cin : out STD_LOGIC;
			sels2 : out STD_LOGIC;
			seldato : out STD_LOGIC;
			selsrc : out STD_LOGIC_VECTOR (2 downto 0);
			seldir : out STD_LOGIC_VECTOR(1 downto 0);
			selop : out STD_LOGIC_VECTOR (3 downto 0);
			selresult : out STD_LOGIC_VECTOR (1 downto 0);
			selc : out STD_LOGIC;
			cadj : out STD_LOGIC;
			selfalgs : out STD_LOGIC_VECTOR (3 downto 0);
			selbranch : out STD_LOGIC_VECTOR (2 downto 0);
			vf : out STD_LOGIC;
			selregw : out STD_LOGIC_VECTOR (2 downto 0);
			memw : out STD_LOGIC;
			seldirw : out STD_LOGIC_VECTOR (1 downto 0));
end u_control;

architecture Behavioral of u_control is
begin
	process (inst)
	begin	
		case inst is
			when X"00C6" => -- LDAB (IMM)
				selregr <= "0000";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '0';
				seldato <= '1';
				selsrc <= "011";
				seldir <= "00";
				selop <= "0100";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf <= '1';
				selregw <= "100";
				memw <= '0';
				seldirw  <= "00";
			when X"0086" => -- LDAA (IMM)
				selregr <= "0000";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '0';
				seldato <= '1';
				selsrc <= "011";
				seldir <= "00";
				selop <= "0100";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf <= '1';
				selregw <= "001";
				memw <= '0';
				seldirw  <= "00";
			when X"001B" => -- ABA (INH)
				selregr <= "0001";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '0';
				seldato <= '0';
				selsrc <= "001";
				seldir <= "00";
				selop <= "0001";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0010";
				selbranch <= "000";
				vf <= '1';
				selregw <= "001";
				memw <= '0';
				seldirw  <= "00";
			when X"007E" => -- JMP (EXT)
				selregr <= "0000";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '0';
				seldato <= '1';
				selsrc <= "011";
				seldir <= "00";
				selop <= "0100";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0000";
				selbranch <= "000";
				vf <= '0';
				selregw <= "000";
				memw <= '0';
				seldirw  <= "00";
			when X"0027" => -- BEQ (REL)
				selregr <= "0000";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '1';
				seldato <= '0';
				selsrc <= "101";
				seldir <= "00";
				selop <= "0001";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0000";
				selbranch <= "010";
				vf <= '1';
				selregw <= "000";
				memw <= '0';
				seldirw  <= "00"; 
			when X"0025" => -- BLO (REL)
				selregr <= "0000";
				sels1 <= '0';
				sr <= '1';
				cin <= '0';
				sels2 <= '1';
				seldato <= '0';
				selsrc <= "101";
				seldir <= "00";
				selop <= "0001";
				selresult <= "01";
				selc <= '1';
				cadj <= '0';
				selfalgs <= "0000";
				selbranch <= "001";
				vf <= '1';
				selregw <= "000";
				memw <= '0';
				seldirw  <= "00";
			when X"0023" => -- BLS (REL)
				selregr  <= "0000";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '1';
				seldato     <= '0';
				selsrc 	  <= "101";
				seldir     <= "00";
				selop 	 <= "0001";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0000";
				selbranch <= "101";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '0';
        seldirw    <= "00";
      when X"0020" => -- BRA (REL)
				selregr  <= "0000";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '1';
				seldato     <= '0';
				selsrc 	  <= "101";
				seldir     <= "00";
				selop 	 <= "0001";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0000";
				selbranch <= "000";
				vf          <= '0';
				selregw   <= "000";
				memw        <= '0';
				seldirw    <= "00";
      when X"007F" => -- CLR (EXT)
				selregr  <= "0000";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '1';
				selsrc 	  <= "010";
				seldir     <= "01";
				selop 	 <= "0011";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0011";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '1';
				seldirw    <= "10";
      when X"0081" => -- CMPA (IMM)
				selregr  <= "0100";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '1';
				selsrc 	  <= "011";
				seldir     <= "01";
				selop 	 <= "0010";
				selresult  <= "00";
				selc        <= '1';
				cadj        <= '1';
				selfalgs <= "0011";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '0';
				seldirw    <= "00";
      when X"00A1" => -- CMPA (IND,X)
				selregr  <= "0110";
				sels1 	    <= '1';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '1';
				selsrc 	  <= "010";
				seldir     <= "00";
				selop 	 <= "0010";
				selresult  <= "00";
				selc        <= '1';
				cadj        <= '1';
				selfalgs <= "0011";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '0';
				seldirw    <= "00";
      when X"007C" => -- INC (EXT)
				selregr  <= "0000";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "010";
				seldir     <= "01";
				selop 	 <= "0001";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '1';
				selfalgs <= "1100";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '1';
				seldirw    <= "10";
      when X"0008" => -- INX (INH)
				selregr  <= "1001";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '1';
				selsrc 	  <= "001";
				seldir     <= "00";
				selop 	 <= "0001";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '1';
				selfalgs <= "0100";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "010";
				memw        <= '0';
				seldirw    <= "00";
      when X"00B6" => -- LDAA (EXT)
				selregr  <= "0000";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "010";
				seldir     <= "01";
				selop 	 <= "0100";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "001";
				memw        <= '0';
				seldirw    <= "00";
      when X"00A6" => -- LDAA (IND,X)
				selregr  <= "1001";
				sels1 	    <= '1';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "010";
				seldir     <= "00";
				selop 	 <= "0100";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "001";
				memw        <= '0';
				seldirw    <= "00";
      when X"00E6" => -- LDAB (IND,X)
				selregr  <= "1001";
				sels1 	    <= '1';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "010";
				seldir     <= "00";
				selop 	 <= "0100";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "100";
				memw        <= '0';
				seldirw    <= "00";
      when X"00CE" => -- LDX (IMM)
				selregr  <= "1001";
				sels1 	    <= '0';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '1';
				selsrc 	  <= "011";
				seldir     <= "00";
				selop 	 <= "0100";
				selresult  <= "01";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "010";
				memw        <= '0';
				seldirw    <= "00";
      when X"00A7" => -- STAA (IND,X)
				selregr  <= "0110";
				sels1 	    <= '1';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "001";
				seldir     <= "00";
				selop 	 <= "0000";
				selresult  <= "11";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '1';
				seldirw    <= "10";
      when X"00E7" => -- STAB (IND,X)
				selregr  <= "0010";
				sels1 	    <= '1';
				sr 			    <= '1';
				cin 		    <= '0';
				sels2 	    <= '0';
				seldato     <= '0';
				selsrc 	  <= "011";
				seldir     <= "00";
				selop 	 <= "0000";
				selresult  <= "11";
				selc        <= '1';
				cadj        <= '0';
				selfalgs <= "0001";
				selbranch <= "000";
				vf          <= '1';
				selregw   <= "000";
				memw        <= '1';
				seldirw    <= "10";
			when others => -- NOP
				selregr <= "0000";
				sels1 <= '0';
				sr <= '0';
				cin <= '0';
				sels2 <= '0';
				seldato <= '0';
				selsrc <= "000";
				seldir <= "00";
				selop <= "0000";
				selresult <= "00";
				selc <= '0';
				cadj <= '0';
				selfalgs <= "0000";
				selbranch <= "000";
				vf <= '1';
				selregw <= "000";
				memw <= '0';
				seldirw  <= "00";				
		end case;
	end process;
end Behavioral;
